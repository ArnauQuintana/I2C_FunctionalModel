module test_I2C();
  
  tb_I2C tb_I2C();
  
  initial
  begin 
     
  #110000 $finish();
  end
  
endmodule
