library verilog;
use verilog.vl_types.all;
entity test_I2C is
end test_I2C;
