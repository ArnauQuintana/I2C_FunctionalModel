library verilog;
use verilog.vl_types.all;
entity tb_I2C is
end tb_I2C;
