library verilog;
use verilog.vl_types.all;
entity sys_rst_fm is
    port(
        Rst_n           : out    vl_logic
    );
end sys_rst_fm;
