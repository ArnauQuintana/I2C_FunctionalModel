library verilog;
use verilog.vl_types.all;
entity sys_clk50MHz_fm is
    port(
        Clk             : out    vl_logic
    );
end sys_clk50MHz_fm;
